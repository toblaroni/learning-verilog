module top #()
(
    input clk,
    output led 
);
endmodule

// Create instance of blinker to pass into top

